module InstructionMem (
    input [31:0] addr,
    output reg [31:0] instruction
);
    parameter ROM_SIZE = 128;
    parameter ROM_BIT  = 7;  // 2^7 = 128
    //reg [31:0] ROM[31:0];

    always @ (*)
        case (addr[ROM_BIT+1:2])
            7'd0: instruction = 32'h08000003;
            7'd1: instruction = 32'h0800004b;
            7'd2: instruction = 32'h08000002;
            7'd3: instruction = 32'h20080014;
            7'd4: instruction = 32'h01000008;
            7'd5: instruction = 32'h3c104000;
            7'd6: instruction = 32'h200bf000;
            7'd7: instruction = 32'hae000008;
            7'd8: instruction = 32'hae0b0000;
            7'd9: instruction = 32'h200cffff;
            7'd10: instruction = 32'h20110000;
            7'd11: instruction = 32'h20120100;
            7'd12: instruction = 32'hae0c0004;
            7'd13: instruction = 32'hae000020;
            7'd14: instruction = 32'h20130000;
            7'd15: instruction = 32'h20080040;
            7'd16: instruction = 32'hae680000;
            7'd17: instruction = 32'h20080079;
            7'd18: instruction = 32'hae680004;
            7'd19: instruction = 32'h20080024;
            7'd20: instruction = 32'hae680008;
            7'd21: instruction = 32'h20080030;
            7'd22: instruction = 32'hae68000c;
            7'd23: instruction = 32'h20080019;
            7'd24: instruction = 32'hae680010;
            7'd25: instruction = 32'h20080012;
            7'd26: instruction = 32'hae680014;
            7'd27: instruction = 32'h20080002;
            7'd28: instruction = 32'hae680018;
            7'd29: instruction = 32'h20080078;
            7'd30: instruction = 32'hae68001c;
            7'd31: instruction = 32'h20080000;
            7'd32: instruction = 32'hae680020;
            7'd33: instruction = 32'h20080010;
            7'd34: instruction = 32'hae680024;
            7'd35: instruction = 32'h20080008;
            7'd36: instruction = 32'hae680028;
            7'd37: instruction = 32'h20080003;
            7'd38: instruction = 32'hae68002c;
            7'd39: instruction = 32'h20080046;
            7'd40: instruction = 32'hae680030;
            7'd41: instruction = 32'h20080021;
            7'd42: instruction = 32'hae680034;
            7'd43: instruction = 32'h20080006;
            7'd44: instruction = 32'hae680038;
            7'd45: instruction = 32'h2008000e;
            7'd46: instruction = 32'hae68003c;
            7'd47: instruction = 32'h8e0e0020;
            7'd48: instruction = 32'h31ce0008;
            7'd49: instruction = 32'h11c0fffd;
            7'd50: instruction = 32'h8e09001c;
            7'd51: instruction = 32'h8e0e0020;
            7'd52: instruction = 32'h31ce0008;
            7'd53: instruction = 32'h11c0fffd;
            7'd54: instruction = 32'h8e0a001c;
            7'd55: instruction = 32'h200d0003;
            7'd56: instruction = 32'h312900ff;
            7'd57: instruction = 32'h314a00ff;
            7'd58: instruction = 32'h00092020;
            7'd59: instruction = 32'h000a2820;
            7'd60: instruction = 32'hae0d0008;
            7'd61: instruction = 32'h112a0007;
            7'd62: instruction = 32'h012a702a;
            7'd63: instruction = 32'h11c00001;
            7'd64: instruction = 32'h08000043;
            7'd65: instruction = 32'h012a4822;
            7'd66: instruction = 32'h0800003d;
            7'd67: instruction = 32'h01495022;
            7'd68: instruction = 32'h0800003d;
            7'd69: instruction = 32'hae090018;
            7'd70: instruction = 32'h8e0e0020;
            7'd71: instruction = 32'h31ce0004;
            7'd72: instruction = 32'h11c0fffd;
            7'd73: instruction = 32'hae09000c;
            7'd74: instruction = 32'h0800002f;
            7'd75: instruction = 32'h8e0d0008;
            7'd76: instruction = 32'h2018fff9;
            7'd77: instruction = 32'h01b86824;
            7'd78: instruction = 32'hae0d0008;
            7'd79: instruction = 32'h12200006;
            7'd80: instruction = 32'h2236ffff;
            7'd81: instruction = 32'h12c00008;
            7'd82: instruction = 32'h22d6ffff;
            7'd83: instruction = 32'h12c0000a;
            7'd84: instruction = 32'h22d6ffff;
            7'd85: instruction = 32'h12c0000c;
            7'd86: instruction = 32'h3088000f;
            7'd87: instruction = 32'h00084080;
            7'd88: instruction = 32'h0113a020;
            7'd89: instruction = 32'h08000066;
            7'd90: instruction = 32'h308800f0;
            7'd91: instruction = 32'h00084082;
            7'd92: instruction = 32'h0113a020;
            7'd93: instruction = 32'h08000066;
            7'd94: instruction = 32'h30a8000f;
            7'd95: instruction = 32'h00084080;
            7'd96: instruction = 32'h0113a020;
            7'd97: instruction = 32'h08000066;
            7'd98: instruction = 32'h30a800f0;
            7'd99: instruction = 32'h00084082;
            7'd100: instruction = 32'h0113a020;
            7'd101: instruction = 32'h08000066;
            7'd102: instruction = 32'h8e950000;
            7'd103: instruction = 32'h02b2a820;
            7'd104: instruction = 32'hae150014;
            7'd105: instruction = 32'h22310001;
            7'd106: instruction = 32'h20080004;
            7'd107: instruction = 32'h12280002;
            7'd108: instruction = 32'h00129040;
            7'd109: instruction = 32'h08000070;
            7'd110: instruction = 32'h20110000;
            7'd111: instruction = 32'h20120100;
            7'd112: instruction = 32'h8e0d0008;
            7'd113: instruction = 32'h35ad0002;
            7'd114: instruction = 32'hae0d0008;
            7'd115: instruction = 32'h03400008;
            default: instruction =32'h8000_0000;
        endcase
endmodule
